library verilog;
use verilog.vl_types.all;
entity CRA_wordslice_vlg_vec_tst is
end CRA_wordslice_vlg_vec_tst;
