library verilog;
use verilog.vl_types.all;
entity PPgen_9bits_vlg_vec_tst is
end PPgen_9bits_vlg_vec_tst;
