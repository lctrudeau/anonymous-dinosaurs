library verilog;
use verilog.vl_types.all;
entity \wordlib8__mbe_1x\ is
    port(
        x0              : in     vl_logic;
        x1              : in     vl_logic;
        x2              : in     vl_logic;
        double          : out    vl_logic;
        neg             : out    vl_logic;
        single          : out    vl_logic;
        vdd             : in     vl_logic;
        gnd             : in     vl_logic
    );
end \wordlib8__mbe_1x\;
