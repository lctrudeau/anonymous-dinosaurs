library verilog;
use verilog.vl_types.all;
entity PosNegUH_sv_unit is
end PosNegUH_sv_unit;
