library verilog;
use verilog.vl_types.all;
entity \wordlib8__PPGen_9bits\ is
    port(
        Double          : in     vl_logic;
        Negate          : in     vl_logic;
        Single          : in     vl_logic;
        Y               : in     vl_logic_vector(0 downto 0);
        Y_1             : in     vl_logic_vector(1 downto 1);
        Y_2             : in     vl_logic_vector(2 downto 2);
        Y_3             : in     vl_logic_vector(3 downto 3);
        Y_4             : in     vl_logic_vector(4 downto 4);
        Y_5             : in     vl_logic_vector(5 downto 5);
        Y_6             : in     vl_logic_vector(6 downto 6);
        Y_7             : in     vl_logic_vector(7 downto 7);
        PP              : out    vl_logic_vector(0 downto 0);
        PP_1            : out    vl_logic_vector(1 downto 1);
        PP_2            : out    vl_logic_vector(2 downto 2);
        PP_3            : out    vl_logic_vector(3 downto 3);
        PP_4            : out    vl_logic_vector(4 downto 4);
        PP_5            : out    vl_logic_vector(5 downto 5);
        PP_6            : out    vl_logic_vector(6 downto 6);
        PP_7            : out    vl_logic_vector(7 downto 7);
        PP_8            : out    vl_logic_vector(8 downto 8);
        Sign            : out    vl_logic;
        vdd             : in     vl_logic;
        vdd_1           : in     vl_logic;
        vdd_1_1         : in     vl_logic;
        vdd_2           : in     vl_logic;
        vdd_3           : in     vl_logic;
        vdd_4           : in     vl_logic;
        vdd_5           : in     vl_logic;
        vdd_6           : in     vl_logic;
        vdd_7           : in     vl_logic;
        vdd_8           : in     vl_logic;
        gnd             : in     vl_logic;
        gnd_1           : in     vl_logic;
        gnd_1_1         : in     vl_logic;
        gnd_2           : in     vl_logic;
        gnd_3           : in     vl_logic;
        gnd_4           : in     vl_logic;
        gnd_5           : in     vl_logic;
        gnd_6           : in     vl_logic;
        gnd_7           : in     vl_logic;
        gnd_8           : in     vl_logic
    );
end \wordlib8__PPGen_9bits\;
