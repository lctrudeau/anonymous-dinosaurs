library verilog;
use verilog.vl_types.all;
entity PosPosLH_sv_unit is
end PosPosLH_sv_unit;
