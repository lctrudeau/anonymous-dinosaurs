library verilog;
use verilog.vl_types.all;
entity PosPosUH_sv_unit is
end PosPosUH_sv_unit;
