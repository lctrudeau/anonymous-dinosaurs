library verilog;
use verilog.vl_types.all;
entity PosZeroLH_sv_unit is
end PosZeroLH_sv_unit;
