// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// PROGRAM		"Quartus II 64-Bit"
// VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"
// CREATED		"Wed Nov 06 13:53:45 2013"

module NAND8_reducer(
	InY,
	Reduced_NAND
);


input wire	[7:0] InY;
output wire	Reduced_NAND;

wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_3;
wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_5;
wire	SYNTHESIZED_WIRE_6;




assign	SYNTHESIZED_WIRE_5 = ~(InY[4] | InY[5]);

assign	SYNTHESIZED_WIRE_4 = ~(InY[2] | InY[3]);

assign	SYNTHESIZED_WIRE_2 =  ~InY[7];

assign	SYNTHESIZED_WIRE_3 = ~(InY[0] | InY[1]);

assign	Reduced_NAND = ~(SYNTHESIZED_WIRE_0 | SYNTHESIZED_WIRE_1);

assign	SYNTHESIZED_WIRE_6 = ~(InY[6] | SYNTHESIZED_WIRE_2);

assign	SYNTHESIZED_WIRE_0 = ~(SYNTHESIZED_WIRE_3 & SYNTHESIZED_WIRE_4);

assign	SYNTHESIZED_WIRE_1 = ~(SYNTHESIZED_WIRE_5 & SYNTHESIZED_WIRE_6);


endmodule
