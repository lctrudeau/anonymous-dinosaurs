library verilog;
use verilog.vl_types.all;
entity NegNegUH_sv_unit is
end NegNegUH_sv_unit;
