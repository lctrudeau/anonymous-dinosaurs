library verilog;
use verilog.vl_types.all;
entity PosNegLH_sv_unit is
end PosNegLH_sv_unit;
