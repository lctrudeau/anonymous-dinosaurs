library verilog;
use verilog.vl_types.all;
entity MBE_vlg_vec_tst is
end MBE_vlg_vec_tst;
