library verilog;
use verilog.vl_types.all;
entity NegNegLH_sv_unit is
end NegNegLH_sv_unit;
