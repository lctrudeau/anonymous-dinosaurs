library verilog;
use verilog.vl_types.all;
entity PosZeroUH_sv_unit is
end PosZeroUH_sv_unit;
