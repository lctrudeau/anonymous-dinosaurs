library verilog;
use verilog.vl_types.all;
entity DUT_vlg_vec_tst is
end DUT_vlg_vec_tst;
