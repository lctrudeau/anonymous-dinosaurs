library verilog;
use verilog.vl_types.all;
entity \wordlib8__PPR\ is
    port(
        PP0             : in     vl_logic_vector(2 downto 2);
        PP0_1           : in     vl_logic_vector(3 downto 3);
        PP0_2           : in     vl_logic_vector(4 downto 4);
        PP0_3           : in     vl_logic_vector(5 downto 5);
        PP0_4           : in     vl_logic_vector(6 downto 6);
        PP0_5           : in     vl_logic_vector(7 downto 7);
        PP0_6           : in     vl_logic_vector(8 downto 8);
        PP1             : in     vl_logic_vector(0 downto 0);
        PP1_1           : in     vl_logic_vector(1 downto 1);
        PP1_2           : in     vl_logic_vector(2 downto 2);
        PP1_3           : in     vl_logic_vector(3 downto 3);
        PP1_4           : in     vl_logic_vector(4 downto 4);
        PP1_5           : in     vl_logic_vector(5 downto 5);
        PP1_6           : in     vl_logic_vector(6 downto 6);
        PP1_7           : in     vl_logic_vector(7 downto 7);
        PP1_8           : in     vl_logic_vector(8 downto 8);
        PP2             : in     vl_logic_vector(0 downto 0);
        PP2_1           : in     vl_logic_vector(1 downto 1);
        PP2_2           : in     vl_logic_vector(2 downto 2);
        PP2_3           : in     vl_logic_vector(3 downto 3);
        PP2_4           : in     vl_logic_vector(4 downto 4);
        PP2_5           : in     vl_logic_vector(5 downto 5);
        PP2_6           : in     vl_logic_vector(6 downto 6);
        PP2_7           : in     vl_logic_vector(7 downto 7);
        PP2_8           : in     vl_logic_vector(8 downto 8);
        PP3             : in     vl_logic_vector(0 downto 0);
        PP3_1           : in     vl_logic_vector(1 downto 1);
        PP3_2           : in     vl_logic_vector(2 downto 2);
        PP3_3           : in     vl_logic_vector(3 downto 3);
        PP3_4           : in     vl_logic_vector(4 downto 4);
        PP3_5           : in     vl_logic_vector(5 downto 5);
        PP3_6           : in     vl_logic_vector(6 downto 6);
        PP3_7           : in     vl_logic_vector(7 downto 7);
        PP3_8           : in     vl_logic_vector(8 downto 8);
        Sign0           : in     vl_logic;
        Sign1           : in     vl_logic;
        Sign2           : in     vl_logic;
        Sign3           : in     vl_logic;
        C0              : out    vl_logic;
        C1              : out    vl_logic;
        C10             : out    vl_logic;
        C11             : out    vl_logic;
        C12             : out    vl_logic;
        C13             : out    vl_logic;
        C2              : out    vl_logic;
        C3              : out    vl_logic;
        C4              : out    vl_logic;
        C5              : out    vl_logic;
        C6              : out    vl_logic;
        C7              : out    vl_logic;
        C8              : out    vl_logic;
        C9              : out    vl_logic;
        S0              : out    vl_logic;
        S1              : out    vl_logic;
        S10             : out    vl_logic;
        S11             : out    vl_logic;
        S12             : out    vl_logic;
        S13             : out    vl_logic;
        S2              : out    vl_logic;
        S3              : out    vl_logic;
        S4              : out    vl_logic;
        S5              : out    vl_logic;
        S6              : out    vl_logic;
        S7              : out    vl_logic;
        S8              : out    vl_logic;
        S9              : out    vl_logic;
        vdd             : in     vl_logic;
        vdd_1           : in     vl_logic;
        vdd_10          : in     vl_logic;
        vdd_11          : in     vl_logic;
        vdd_12          : in     vl_logic;
        vdd_1_1         : in     vl_logic;
        vdd_2           : in     vl_logic;
        vdd_3           : in     vl_logic;
        vdd_4           : in     vl_logic;
        vdd_5           : in     vl_logic;
        vdd_6           : in     vl_logic;
        vdd_7           : in     vl_logic;
        vdd_8           : in     vl_logic;
        vdd_9           : in     vl_logic;
        gnd             : in     vl_logic;
        gnd_1           : in     vl_logic;
        gnd_10          : in     vl_logic;
        gnd_11          : in     vl_logic;
        gnd_12          : in     vl_logic;
        gnd_1_1         : in     vl_logic;
        gnd_2           : in     vl_logic;
        gnd_3           : in     vl_logic;
        gnd_4           : in     vl_logic;
        gnd_5           : in     vl_logic;
        gnd_6           : in     vl_logic;
        gnd_7           : in     vl_logic;
        gnd_8           : in     vl_logic;
        gnd_9           : in     vl_logic
    );
end \wordlib8__PPR\;
