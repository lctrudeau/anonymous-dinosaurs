library verilog;
use verilog.vl_types.all;
entity MBE_wordslice_vlg_vec_tst is
end MBE_wordslice_vlg_vec_tst;
