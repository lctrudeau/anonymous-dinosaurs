library verilog;
use verilog.vl_types.all;
entity \wordlib8__CPA\ is
    port(
        a0              : in     vl_logic;
        a1              : in     vl_logic;
        a10             : in     vl_logic;
        a11             : in     vl_logic;
        a12             : in     vl_logic;
        a13             : in     vl_logic;
        a2              : in     vl_logic;
        a3              : in     vl_logic;
        a4              : in     vl_logic;
        a5              : in     vl_logic;
        a6              : in     vl_logic;
        a7              : in     vl_logic;
        a8              : in     vl_logic;
        a9              : in     vl_logic;
        b0              : in     vl_logic;
        b1              : in     vl_logic;
        b10             : in     vl_logic;
        b11             : in     vl_logic;
        b12             : in     vl_logic;
        b13             : in     vl_logic;
        b2              : in     vl_logic;
        b3              : in     vl_logic;
        b4              : in     vl_logic;
        b5              : in     vl_logic;
        b6              : in     vl_logic;
        b7              : in     vl_logic;
        b8              : in     vl_logic;
        b9              : in     vl_logic;
        cout            : out    vl_logic;
        s0              : out    vl_logic;
        s1              : out    vl_logic;
        s10             : out    vl_logic;
        s11             : out    vl_logic;
        s12             : out    vl_logic;
        s13             : out    vl_logic;
        s2              : out    vl_logic;
        s3              : out    vl_logic;
        s4              : out    vl_logic;
        s5              : out    vl_logic;
        s6              : out    vl_logic;
        s7              : out    vl_logic;
        s8              : out    vl_logic;
        s9              : out    vl_logic;
        vdd             : in     vl_logic;
        vdd_1           : in     vl_logic;
        vdd_10          : in     vl_logic;
        vdd_11          : in     vl_logic;
        vdd_12          : in     vl_logic;
        vdd_1_1         : in     vl_logic;
        vdd_2           : in     vl_logic;
        vdd_3           : in     vl_logic;
        vdd_4           : in     vl_logic;
        vdd_5           : in     vl_logic;
        vdd_6           : in     vl_logic;
        vdd_7           : in     vl_logic;
        vdd_8           : in     vl_logic;
        vdd_9           : in     vl_logic;
        gnd             : in     vl_logic;
        gnd_1           : in     vl_logic;
        gnd_10          : in     vl_logic;
        gnd_11          : in     vl_logic;
        gnd_12          : in     vl_logic;
        gnd_1_1         : in     vl_logic;
        gnd_2           : in     vl_logic;
        gnd_3           : in     vl_logic;
        gnd_4           : in     vl_logic;
        gnd_5           : in     vl_logic;
        gnd_6           : in     vl_logic;
        gnd_7           : in     vl_logic;
        gnd_8           : in     vl_logic;
        gnd_9           : in     vl_logic
    );
end \wordlib8__CPA\;
